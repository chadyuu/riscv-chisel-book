../../../chisel-template/rtl/riscv/top.sv